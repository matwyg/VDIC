/*
asdf
*/